// Author: Ratnodeep Bandyopadhyay. Copyright 2022.
// Simplify Module


module turn_positive


module simplify #(INT_WIDTH = 64, THRESH_INDEX = 30)
    (
        input [INT_WIDTH-1:0] in_num,
        input [INT_WIDTH-1:0] in_den,
        input clk,

        output [INT_WIDTH-2:0] out_num,
        output [INT_WIDTH-1:0] out_den
    )

    reg

    

    always @(posedge clk) begin
        

    end

endmodule
